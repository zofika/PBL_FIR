////////////////////////////////////////////////////////////////////////
//   główny moduł dla FIR.
//   Do testów w cocoTB
///////////////////////////////////////////////////////////////////////


//FSM

//Licznik

//Licznik petli  

//Shift R

//Acc

//sumator

//mnozenie
