////////////////////////////////////////////////////////////////////////
//   główny moduł dla APB.
//   Do testów w cocoTB
///////////////////////////////////////////////////////////////////////



//APB

//CDC

//Dekoder

//MUX'y
//MUX_DEKODER

//MUX_CDC_wsp

//RAM (tutaj jest jeszcze ten AND - ale może bez niego?)

//Rejestry sterujace
