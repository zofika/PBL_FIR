////////////////////////////////////////////////////////////////////////
//   główny moduł dla AXI.
//   Do testów w cocoTB
///////////////////////////////////////////////////////////////////////

//AXI


//MUX'y


//RAM (wej)


//RAM (wyj)
