////////////////////////////////////////////////////////////////////////
//   główny moduł dla APB.
//   Do testów w cocoTB
///////////////////////////////////////////////////////////////////////



//APB


//CDC


//Dekoder

//MUX'y

//RAM

//Rejestry sterujace

