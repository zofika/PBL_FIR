////////////////////////////////////////////////////////////////////////
//   główny moduł dla naszego projektu.
///////////////////////////////////////////////////////////////////////


//APB_main


//AXI_main


//FIR_main


